
module clock (
	clk_clk,
	clk_25m_clk,
	clk_116800_clk,
	clk_12m_clk,
	reset_reset_n);	

	input		clk_clk;
	output		clk_25m_clk;
	output		clk_116800_clk;
	output		clk_12m_clk;
	input		reset_reset_n;
endmodule
